LIBRARY ieee;
CONTEXT ieee.ieee_std_context;

USE work.RiscVPkg.ALL;

ENTITY Cpu IS
    PORT (
        clk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        halt : OUT STD_LOGIC := '0'
    );
END ENTITY Cpu;

ARCHITECTURE rtl OF Cpu IS
    SIGNAL pc : STD_LOGIC_VECTOR(XLEN - 1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL registerFile : RegistersType;

    SIGNAL rs1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
    SIGNAL rs2 : STD_LOGIC_VECTOR(4 DOWNTO 0);
    SIGNAL rd : STD_LOGIC_VECTOR(4 DOWNTO 0);
    SIGNAL immediate : STD_LOGIC_VECTOR(31 DOWNTO 0);

    SIGNAL instType : InstructionType;
    SIGNAL instruction : STD_LOGIC_VECTOR(31 DOWNTO 0);

    SIGNAL wr_addr : STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
    SIGNAL wr_data : STD_LOGIC_VECTOR(XLEN - 1 DOWNTO 0);
    SIGNAL wr_strobe : STD_LOGIC;

    SIGNAL ram_we : STD_LOGIC;
    SIGNAL ram_di : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL ram_do : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL ram_addr : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
BEGIN
    -- halt once we hit an ebreak
    halt <= '1' WHEN instType = EBREAK ELSE
        '0';

    PROCESS (clk)
    BEGIN
        IF rising_edge(clk) THEN
            IF reset = '1' THEN
                pc <= (OTHERS => '0');
            ELSE
                pc <= STD_LOGIC_VECTOR(UNSIGNED(pc) + 4);
            END IF;
        END IF;
    END PROCESS;

    -- temp ram instruction read
    instruction <= ram_do;
    ram_addr <= pc;

    Registers_inst : ENTITY work.Registers
        PORT MAP(
            clk => clk,
            reset => reset,
            --pc => pc,
            registersValue => registerFile,
            wr_addr => to_integer(unsigned(wr_addr)),
            wr_data => wr_data,
            wr_strobe => wr_strobe
        );

    Ram_inst : ENTITY work.Ram
        PORT MAP(
            clk => clk,
            we => ram_we,
            -- word-addressed
            addr => ram_addr(7 DOWNTO 2),
            di => ram_di,
            do => ram_do
        );

    InstructionDecoder_inst : ENTITY work.InstructionDecoder
        PORT MAP(
            instructionType => instType,
            instruction => instruction,
            immediate => immediate,
            rs1 => rs1,
            rs2 => rs2,
            rd => rd
        );
END ARCHITECTURE;